// --------------------------------------------------------------------------------------------------------------------
// IP Block    : MESH
// Function    : Network
// Module name : MESH_Network
// Description : Instantiates a 2D Mesh Network of routers
// Uses        : MESH_Router.sv
// Notes       : Incomplete
// --------------------------------------------------------------------------------------------------------------------

`include "config.sv"

module MESH_network