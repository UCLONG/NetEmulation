// IP Block    : MESH
// Sub Block   :
// Function    :
// Module name :
// Description :
// Uses        :
// Notes       :

`include "config.sv"

