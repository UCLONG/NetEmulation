// `define VC