// IP Block    : SO
// Function    : Network
// Module name : SO_Network
// Description :
// Uses        : config.sv, SO_AllocSimple.sv, SO_TxSimple.sv and SO_PhotonicSwitch.sv
// Notes       :
