module FIFO
 
  // The width and the depth of the FIFO is paramatised.  Standard set as a 4 deep 64 bit memory.
 
  #(parameter FIFO_WIDTH = 64,
    parameter FIFO_DEPTH = 4)
   
   (output reg    [FIFO_WIDTH-1:0] dataOut,
    output logic  full, empty, write_ack, read_valid,
     
     input reg    [FIFO_WIDTH-1:0] dataIn, 
     input logic  read, write, clk);
     
     
  // Function to calculate Log2(n)
  
  function int log2
    (input int n);
    
    begin
      log2 = 0;     // log2 is zero to start
      n--;          // decrement 'n'
      while (n > 0) // While n is greater than 0
        begin
          log2++;   // Increment 'log2'
          n >>= 1;  // Bitwise shift 'n' to the right by one position
        end
    end
    
  endfunction
  
  
  // Declare Memory Array of 'MEM_DEPTH', 'MEM_WIDTH' bit words.
  // Default Memory Array of 4, 64 bit words.
  
  reg [FIFO_WIDTH-1:0] FIFO [0:FIFO_DEPTH-1];
  
  
  // Control Flags (read_ptr, write_ptr, full, empty).  The read and write pointers are calculated using a binary representation for each cell.
  // Each pointer has one more significant bit than required.  This enables comparison to check if the FIFO is full or empty. 
  
  reg [log2(MEM_DEPTH):0] read_ptr, write_ptr;  // Note the inclusion of an extra significant bit.
  assign empty = (write_ptr == read_ptr);       // If the write and read pointers including their MSB are equal, the FIFO is empty.
  assign full  = ((write_ptr[log2(FIFO_DEPTH)-1:0] == read_ptr[log2(FIFO_DEPTH)-1:0]) && write_ptr[Log2(FIFO_DEPTH)] ^ read_ptr[log2(FIFO_DEPTH)]);
  
  
  // Memory Read and Write on the rising edge of the clock, with write acknowledgement.
  
  always_ff @ (posedge clk)
    begin
      if (read && ~empty)                             // If the read signal is asserted and the FIFO is not empty
        begin
        dataOut <= mem[read_ptr[log2(MEM_DEPTH)-1]];  // dataOut will be read from the memory
        read_valid <= 1'b0;                           // A Valid signal will be asserted to indicate the data on dataOut is valid
        read_ptr++;                                   // The read_ptr is incremented, truncating if to big.
        end
      if (write && ~full)                             // If the write signal is asserted and the FIFO is not full
        begin                             
        mem[write_ptr[log2(MEM_DEPTH)-1]] <= dataIn;  // dataIn will be written to memory
        write_ack <= 1'b1;                            // A write acknowledgement signal will be asserted to indicate write has worked
        write_ptr++;                                  // The write pointer is incremented, truncating if to big.
        end
      else                                            // Otherwise
        write_ack <= 1'b0;                            // The write is not acknowledged
        read_valid <= 1'b0;                           // The read date is not valid
    end

endmodule