// `define VC
// `define iSLIP

`define MESH
// `define TORUS