// `define VC
// `define iSLIP
// `define TORUS